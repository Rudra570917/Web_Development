<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>3.55271e-015,-1.42109e-014,122.4,-60.5</PageViewport>
<gate>
<ID>2</ID>
<type>BE_JKFF_LOW_NT</type>
<position>38,-28.5</position>
<input>
<ID>J</ID>1 </input>
<input>
<ID>K</ID>1 </input>
<output>
<ID>Q</ID>4 </output>
<input>
<ID>clock</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>4</ID>
<type>BE_JKFF_LOW_NT</type>
<position>52.5,-28.5</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>5 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>23,-23</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>BB_CLOCK</type>
<position>21.5,-29</position>
<output>
<ID>CLK</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>10</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>62,-29</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>40.5,-19</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-30.5,32,-23.5</points>
<intersection>-30.5 2</intersection>
<intersection>-26.5 1</intersection>
<intersection>-23.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-26.5,35,-26.5</points>
<connection>
<GID>2</GID>
<name>J</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-30.5,35,-30.5</points>
<connection>
<GID>2</GID>
<name>K</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>28,-23.5,32,-23.5</points>
<intersection>28 5</intersection>
<intersection>32 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>28,-23.5,28,-23</points>
<intersection>-23.5 4</intersection>
<intersection>-23 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>25,-23,28,-23</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>28 5</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-31.5,48,-25.5</points>
<intersection>-31.5 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-25.5,48.5,-25.5</points>
<intersection>48 0</intersection>
<intersection>48.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-31.5,49.5,-31.5</points>
<intersection>48 0</intersection>
<intersection>49.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48.5,-25.5,48.5,-25</points>
<intersection>-25.5 1</intersection>
<intersection>-25 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-25,48.5,-25</points>
<intersection>42.5 8</intersection>
<intersection>43.5 5</intersection>
<intersection>48.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>43.5,-26.5,43.5,-25</points>
<intersection>-26.5 6</intersection>
<intersection>-25 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>43.5,-26.5,49.5,-26.5</points>
<connection>
<GID>4</GID>
<name>J</name></connection>
<intersection>43.5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>49.5,-31.5,49.5,-30.5</points>
<connection>
<GID>4</GID>
<name>K</name></connection>
<intersection>-31.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>42.5,-25,42.5,-19</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-25 4</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-29,30,-28.5</points>
<intersection>-29 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-28.5,35,-28.5</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-29,30,-29</points>
<connection>
<GID>8</GID>
<name>CLK</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-28.5,45,-27.5</points>
<intersection>-28.5 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-28.5,59,-28.5</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>45 0</intersection>
<intersection>59 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-27.5,45,-27.5</points>
<intersection>41 3</intersection>
<intersection>45 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41,-27.5,41,-26.5</points>
<connection>
<GID>2</GID>
<name>Q</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>59,-30,59,-28.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-29,57,-26.5</points>
<intersection>-29 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-29,59,-29</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-26.5,57,-26.5</points>
<connection>
<GID>4</GID>
<name>Q</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>