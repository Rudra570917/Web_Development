<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>5.1981,21.9113,295.659,-121.658</PageViewport>
<gate>
<ID>4</ID>
<type>BE_JKFF_LOW</type>
<position>34,-27</position>
<input>
<ID>J</ID>5 </input>
<input>
<ID>K</ID>5 </input>
<output>
<ID>Q</ID>3 </output>
<input>
<ID>clear</ID>8 </input>
<input>
<ID>clock</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5</ID>
<type>BE_JKFF_LOW</type>
<position>44,-27</position>
<input>
<ID>J</ID>5 </input>
<input>
<ID>K</ID>5 </input>
<output>
<ID>Q</ID>4 </output>
<input>
<ID>clear</ID>8 </input>
<input>
<ID>clock</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>BE_JKFF_LOW</type>
<position>54,-27</position>
<input>
<ID>J</ID>5 </input>
<input>
<ID>K</ID>5 </input>
<output>
<ID>Q</ID>6 </output>
<input>
<ID>clear</ID>8 </input>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7</ID>
<type>BE_JKFF_LOW</type>
<position>64,-27</position>
<input>
<ID>J</ID>5 </input>
<input>
<ID>K</ID>5 </input>
<output>
<ID>Q</ID>1 </output>
<input>
<ID>clear</ID>8 </input>
<input>
<ID>clock</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>11</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>77,-27</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>1 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>25,-20.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_AND2</type>
<position>203,-20</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>182 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_AND2</type>
<position>203.5,-26</position>
<input>
<ID>IN_0</ID>177 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>BA_NAND2</type>
<position>77,-16.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>AE_OR2</type>
<position>211,-23</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>180 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_AND3</type>
<position>229,-14</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>182 </input>
<input>
<ID>IN_2</ID>185 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>17</ID>
<type>BB_CLOCK</type>
<position>24.5,-27</position>
<output>
<ID>CLK</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_AND3</type>
<position>229,-22</position>
<input>
<ID>IN_0</ID>177 </input>
<input>
<ID>IN_1</ID>183 </input>
<input>
<ID>IN_2</ID>186 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>211</ID>
<type>AE_OR2</type>
<position>236,-18</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>254,-28</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>186 </input>
<input>
<ID>IN_2</ID>190 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>213</ID>
<type>BB_CLOCK</type>
<position>184,-38</position>
<output>
<ID>CLK</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_LABEL</type>
<position>209.5,-8</position>
<gparam>LABEL_TEXT 3 bit Sync Up/Down Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_TOGGLE</type>
<position>186,-19</position>
<output>
<ID>OUT_0</ID>177 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_TOGGLE</type>
<position>186,-25</position>
<output>
<ID>OUT_0</ID>178 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>217</ID>
<type>AE_SMALL_INVERTER</type>
<position>194,-19</position>
<input>
<ID>IN_0</ID>177 </input>
<output>
<ID>OUT_0</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>BE_JKFF_LOW</type>
<position>194,-31</position>
<input>
<ID>J</ID>178 </input>
<input>
<ID>K</ID>178 </input>
<output>
<ID>Q</ID>183 </output>
<input>
<ID>clock</ID>191 </input>
<output>
<ID>nQ</ID>182 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>219</ID>
<type>BE_JKFF_LOW</type>
<position>219,-29</position>
<input>
<ID>J</ID>184 </input>
<input>
<ID>K</ID>184 </input>
<output>
<ID>Q</ID>186 </output>
<input>
<ID>clock</ID>191 </input>
<output>
<ID>nQ</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>220</ID>
<type>BE_JKFF_LOW</type>
<position>244,-29</position>
<input>
<ID>J</ID>189 </input>
<input>
<ID>K</ID>189 </input>
<output>
<ID>Q</ID>190 </output>
<input>
<ID>clock</ID>191 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>49</ID>
<type>BB_CLOCK</type>
<position>31,-51.5</position>
<output>
<ID>CLK</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>24,-43</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_AND2</type>
<position>48,-48.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>48,-54.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_OR2</type>
<position>56.5,-51.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>BE_JKFF_LOW_NT</type>
<position>40,-51.5</position>
<input>
<ID>J</ID>49 </input>
<input>
<ID>K</ID>49 </input>
<output>
<ID>Q</ID>46 </output>
<input>
<ID>clock</ID>42 </input>
<output>
<ID>nQ</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>55</ID>
<type>BE_JKFF_LOW_NT</type>
<position>65,-51.5</position>
<input>
<ID>J</ID>49 </input>
<input>
<ID>K</ID>49 </input>
<output>
<ID>Q</ID>44 </output>
<input>
<ID>clock</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>56</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>74,-52</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>44 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>57</ID>
<type>AE_SMALL_INVERTER</type>
<position>38,-43</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>33,-45.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>71</ID>
<type>BB_CLOCK</type>
<position>31,-80.5</position>
<output>
<ID>CLK</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>26.5,-68</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>48,-77.5</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_AND2</type>
<position>48,-83.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AE_OR2</type>
<position>56.5,-80.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>BE_JKFF_LOW_NT</type>
<position>40,-80.5</position>
<input>
<ID>J</ID>68 </input>
<input>
<ID>K</ID>68 </input>
<output>
<ID>Q</ID>66 </output>
<input>
<ID>clock</ID>63 </input>
<output>
<ID>nQ</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>77</ID>
<type>BE_JKFF_LOW_NT</type>
<position>65,-80.5</position>
<input>
<ID>J</ID>68 </input>
<input>
<ID>K</ID>68 </input>
<output>
<ID>Q</ID>65 </output>
<input>
<ID>clock</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>78</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>74,-78.5</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>65 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_TOGGLE</type>
<position>33,-74.5</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>80</ID>
<type>AE_SMALL_INVERTER</type>
<position>26.5,-76</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>122.5,-8.5</position>
<gparam>LABEL_TEXT 3 bit Sync Up Counter using JK FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>BE_JKFF_LOW</type>
<position>108,-23</position>
<input>
<ID>J</ID>128 </input>
<input>
<ID>K</ID>128 </input>
<output>
<ID>Q</ID>129 </output>
<input>
<ID>clock</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>147</ID>
<type>BE_JKFF_LOW</type>
<position>118,-23</position>
<input>
<ID>J</ID>129 </input>
<input>
<ID>K</ID>129 </input>
<output>
<ID>Q</ID>131 </output>
<input>
<ID>clock</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>148</ID>
<type>BE_JKFF_LOW</type>
<position>134,-23</position>
<input>
<ID>J</ID>130 </input>
<input>
<ID>K</ID>130 </input>
<output>
<ID>Q</ID>132 </output>
<input>
<ID>clock</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_TOGGLE</type>
<position>99,-16</position>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>150</ID>
<type>BB_CLOCK</type>
<position>98,-28</position>
<output>
<ID>CLK</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_AND2</type>
<position>126,-15</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>152</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>143,-22</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>131 </input>
<input>
<ID>IN_2</ID>132 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>124.5,-35.5</position>
<gparam>LABEL_TEXT 3 bit Sync Down Counter using JK FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>BE_JKFF_LOW</type>
<position>108,-50</position>
<input>
<ID>J</ID>134 </input>
<input>
<ID>K</ID>134 </input>
<output>
<ID>Q</ID>140 </output>
<input>
<ID>clock</ID>133 </input>
<output>
<ID>nQ</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>155</ID>
<type>BE_JKFF_LOW</type>
<position>118,-50</position>
<input>
<ID>J</ID>137 </input>
<input>
<ID>K</ID>137 </input>
<output>
<ID>Q</ID>139 </output>
<input>
<ID>clock</ID>133 </input>
<output>
<ID>nQ</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>156</ID>
<type>BE_JKFF_LOW</type>
<position>134,-50</position>
<input>
<ID>J</ID>135 </input>
<input>
<ID>K</ID>135 </input>
<output>
<ID>Q</ID>136 </output>
<input>
<ID>clock</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>99,-43</position>
<output>
<ID>OUT_0</ID>134 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>158</ID>
<type>BB_CLOCK</type>
<position>98,-55</position>
<output>
<ID>CLK</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND2</type>
<position>126,-42</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>143,-49</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>139 </input>
<input>
<ID>IN_2</ID>136 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>125,-60</position>
<gparam>LABEL_TEXT MOD 10 Sync Up Counter using JK FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>BE_JKFF_LOW</type>
<position>107,-77</position>
<input>
<ID>J</ID>142 </input>
<input>
<ID>K</ID>142 </input>
<output>
<ID>Q</ID>147 </output>
<input>
<ID>clock</ID>141 </input>
<output>
<ID>nQ</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>163</ID>
<type>BE_JKFF_LOW</type>
<position>123,-77</position>
<input>
<ID>J</ID>149 </input>
<input>
<ID>K</ID>147 </input>
<output>
<ID>Q</ID>144 </output>
<input>
<ID>clock</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>164</ID>
<type>BE_JKFF_LOW</type>
<position>139,-76.5</position>
<input>
<ID>J</ID>150 </input>
<input>
<ID>K</ID>150 </input>
<output>
<ID>Q</ID>143 </output>
<input>
<ID>clock</ID>141 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_TOGGLE</type>
<position>99,-70</position>
<output>
<ID>OUT_0</ID>142 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>166</ID>
<type>BB_CLOCK</type>
<position>97,-81.5</position>
<output>
<ID>CLK</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_AND2</type>
<position>131,-67.5</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>169,-75.5</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_2</ID>143 </input>
<input>
<ID>IN_3</ID>145 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 9</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>169</ID>
<type>BE_JKFF_LOW</type>
<position>158,-75.5</position>
<input>
<ID>J</ID>151 </input>
<input>
<ID>K</ID>147 </input>
<output>
<ID>Q</ID>145 </output>
<input>
<ID>clock</ID>141 </input>
<output>
<ID>nQ</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND2</type>
<position>115,-67.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_AND3</type>
<position>150,-69.5</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_2</ID>143 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>172</ID>
<type>BE_JKFF_LOW</type>
<position>130,-106</position>
<input>
<ID>J</ID>155 </input>
<input>
<ID>K</ID>155 </input>
<output>
<ID>Q</ID>159 </output>
<input>
<ID>clock</ID>152 </input>
<output>
<ID>nQ</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>173</ID>
<type>BE_JKFF_LOW</type>
<position>146,-106</position>
<input>
<ID>J</ID>161 </input>
<input>
<ID>K</ID>161 </input>
<output>
<ID>Q</ID>158 </output>
<input>
<ID>clock</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>174</ID>
<type>BE_JKFF_LOW</type>
<position>156,-106</position>
<input>
<ID>J</ID>158 </input>
<input>
<ID>K</ID>158 </input>
<output>
<ID>Q</ID>160 </output>
<input>
<ID>clock</ID>152 </input>
<output>
<ID>nQ</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>175</ID>
<type>BB_CLOCK</type>
<position>120,-114.5</position>
<output>
<ID>CLK</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_AND2</type>
<position>115,-96</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_AND2</type>
<position>115,-102</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>AE_OR2</type>
<position>122,-99</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AE_OR2</type>
<position>138.5,-100.5</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>167,-105</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>158 </input>
<input>
<ID>IN_2</ID>160 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67,-25,74,-25</points>
<connection>
<GID>7</GID>
<name>Q</name></connection>
<connection>
<GID>11</GID>
<name>IN_3</name></connection>
<intersection>73 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>73,-25,73,-17.5</points>
<intersection>-25 1</intersection>
<intersection>-17.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>73,-17.5,74,-17.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>73 6</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-35,73,-35</points>
<intersection>38 3</intersection>
<intersection>73 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-35,38,-25</points>
<intersection>-35 1</intersection>
<intersection>-27 8</intersection>
<intersection>-25 7</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>73,-35,73,-28</points>
<intersection>-35 1</intersection>
<intersection>-28 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>73,-28,74,-28</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>73 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>37,-25,38,-25</points>
<connection>
<GID>4</GID>
<name>Q</name></connection>
<intersection>38 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>38,-27,41,-27</points>
<connection>
<GID>5</GID>
<name>clock</name></connection>
<intersection>38 3</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-34,49,-25</points>
<intersection>-34 1</intersection>
<intersection>-27 6</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-34,72,-34</points>
<intersection>49 0</intersection>
<intersection>72 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,-25,49,-25</points>
<connection>
<GID>5</GID>
<name>Q</name></connection>
<intersection>49 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>72,-34,72,-15.5</points>
<intersection>-34 1</intersection>
<intersection>-27 7</intersection>
<intersection>-15.5 13</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>49,-27,51,-27</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>72,-27,74,-27</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>72 4</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>72,-15.5,74,-15.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>72 4</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-20.5,60,-20.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>30 3</intersection>
<intersection>40 6</intersection>
<intersection>50 8</intersection>
<intersection>60 10</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>30,-29,30,-20.5</points>
<intersection>-29 11</intersection>
<intersection>-25 12</intersection>
<intersection>-20.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>40,-29,40,-20.5</points>
<intersection>-29 13</intersection>
<intersection>-25 14</intersection>
<intersection>-20.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>50,-29,50,-20.5</points>
<intersection>-29 15</intersection>
<intersection>-25 16</intersection>
<intersection>-20.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>60,-29,60,-20.5</points>
<intersection>-29 17</intersection>
<intersection>-25 18</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>30,-29,31,-29</points>
<connection>
<GID>4</GID>
<name>K</name></connection>
<intersection>30 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>30,-25,31,-25</points>
<connection>
<GID>4</GID>
<name>J</name></connection>
<intersection>30 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>40,-29,41,-29</points>
<connection>
<GID>5</GID>
<name>K</name></connection>
<intersection>40 6</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>40,-25,41,-25</points>
<connection>
<GID>5</GID>
<name>J</name></connection>
<intersection>40 6</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>50,-29,51,-29</points>
<connection>
<GID>6</GID>
<name>K</name></connection>
<intersection>50 8</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>50,-25,51,-25</points>
<connection>
<GID>6</GID>
<name>J</name></connection>
<intersection>50 8</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>60,-29,61,-29</points>
<connection>
<GID>7</GID>
<name>K</name></connection>
<intersection>60 10</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>60,-25,61,-25</points>
<connection>
<GID>7</GID>
<name>J</name></connection>
<intersection>60 10</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-33,59,-25</points>
<intersection>-33 1</intersection>
<intersection>-27 6</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-33,71,-33</points>
<intersection>59 0</intersection>
<intersection>71 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-25,59,-25</points>
<connection>
<GID>6</GID>
<name>Q</name></connection>
<intersection>59 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-33,71,-26</points>
<intersection>-33 1</intersection>
<intersection>-26 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>71,-26,74,-26</points>
<connection>
<GID>11</GID>
<name>IN_2</name></connection>
<intersection>71 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>59,-27,61,-27</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-27,31,-27</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<connection>
<GID>17</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-32,64,-31</points>
<connection>
<GID>7</GID>
<name>clear</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-32,81,-32</points>
<intersection>34 6</intersection>
<intersection>44 7</intersection>
<intersection>54 8</intersection>
<intersection>64 0</intersection>
<intersection>81 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>81,-32,81,-16.5</points>
<intersection>-32 1</intersection>
<intersection>-16.5 9</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>34,-32,34,-31</points>
<connection>
<GID>4</GID>
<name>clear</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>44,-32,44,-31</points>
<connection>
<GID>5</GID>
<name>clear</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>54,-32,54,-31</points>
<connection>
<GID>6</GID>
<name>clear</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>80,-16.5,81,-16.5</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>81 2</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-50.5,52.5,-48.5</points>
<intersection>-50.5 1</intersection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-50.5,53.5,-50.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-48.5,52.5,-48.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-54.5,52.5,-52.5</points>
<intersection>-54.5 2</intersection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-52.5,53.5,-52.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-54.5,52.5,-54.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-51.5,37,-51.5</points>
<connection>
<GID>49</GID>
<name>CLK</name></connection>
<connection>
<GID>54</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-51.5,62,-51.5</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<connection>
<GID>55</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-52,70,-49.5</points>
<intersection>-52 1</intersection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-52,71,-52</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-49.5,70,-49.5</points>
<connection>
<GID>55</GID>
<name>Q</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-47.5,44,-43</points>
<intersection>-47.5 3</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>40,-43,44,-43</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>44,-47.5,45,-47.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-58.5,70,-58.5</points>
<intersection>44 8</intersection>
<intersection>70 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>70,-58.5,70,-53</points>
<intersection>-58.5 1</intersection>
<intersection>-53 11</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>44,-58.5,44,-49.5</points>
<intersection>-58.5 1</intersection>
<intersection>-49.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>43,-49.5,45,-49.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<connection>
<GID>54</GID>
<name>Q</name></connection>
<intersection>44 8</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>70,-53,71,-53</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>70 7</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>27,-57,27,-43</points>
<intersection>-57 4</intersection>
<intersection>-43 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>27,-57,43,-57</points>
<intersection>27 3</intersection>
<intersection>43 8</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>26,-43,36,-43</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>43,-57,43,-55.5</points>
<intersection>-57 4</intersection>
<intersection>-55.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>43,-55.5,45,-55.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>43 8</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-53.5,45,-53.5</points>
<connection>
<GID>54</GID>
<name>nQ</name></connection>
<connection>
<GID>52</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-53.5,36,-45.5</points>
<intersection>-53.5 4</intersection>
<intersection>-49.5 9</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-45.5,61,-45.5</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection>
<intersection>61 6</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36,-53.5,37,-53.5</points>
<connection>
<GID>54</GID>
<name>K</name></connection>
<intersection>36 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>61,-53.5,61,-45.5</points>
<intersection>-53.5 10</intersection>
<intersection>-49.5 11</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>36,-49.5,37,-49.5</points>
<connection>
<GID>54</GID>
<name>J</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>61,-53.5,62,-53.5</points>
<connection>
<GID>55</GID>
<name>K</name></connection>
<intersection>61 6</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>61,-49.5,62,-49.5</points>
<connection>
<GID>55</GID>
<name>J</name></connection>
<intersection>61 6</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-79.5,52.5,-77.5</points>
<intersection>-79.5 1</intersection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-79.5,53.5,-79.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-77.5,52.5,-77.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-83.5,52.5,-81.5</points>
<intersection>-83.5 2</intersection>
<intersection>-81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-81.5,53.5,-81.5</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-83.5,52.5,-83.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-80.5,37,-80.5</points>
<connection>
<GID>76</GID>
<name>clock</name></connection>
<connection>
<GID>71</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59.5,-80.5,62,-80.5</points>
<connection>
<GID>77</GID>
<name>clock</name></connection>
<connection>
<GID>75</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-78.5,71,-78.5</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<connection>
<GID>77</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-87.5,70,-87.5</points>
<intersection>44 8</intersection>
<intersection>70 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>70,-87.5,70,-79.5</points>
<intersection>-87.5 1</intersection>
<intersection>-79.5 14</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>44,-87.5,44,-78.5</points>
<intersection>-87.5 1</intersection>
<intersection>-78.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>43,-78.5,45,-78.5</points>
<connection>
<GID>76</GID>
<name>Q</name></connection>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>44 8</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>70,-79.5,71,-79.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>70 7</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-82.5,45,-82.5</points>
<connection>
<GID>76</GID>
<name>nQ</name></connection>
<connection>
<GID>74</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-82.5,36,-74.5</points>
<intersection>-82.5 4</intersection>
<intersection>-78.5 9</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-74.5,61,-74.5</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection>
<intersection>61 6</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36,-82.5,37,-82.5</points>
<connection>
<GID>76</GID>
<name>K</name></connection>
<intersection>36 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>61,-82.5,61,-74.5</points>
<intersection>-82.5 10</intersection>
<intersection>-78.5 11</intersection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>36,-78.5,37,-78.5</points>
<connection>
<GID>76</GID>
<name>J</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>61,-82.5,62,-82.5</points>
<connection>
<GID>77</GID>
<name>K</name></connection>
<intersection>61 6</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>61,-78.5,62,-78.5</points>
<connection>
<GID>77</GID>
<name>J</name></connection>
<intersection>61 6</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-74,26.5,-70</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-71.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-71.5,44,-71.5</points>
<intersection>26.5 0</intersection>
<intersection>44 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>44,-76.5,44,-71.5</points>
<intersection>-76.5 8</intersection>
<intersection>-71.5 3</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>44,-76.5,45,-76.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>44 4</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-85.5,26.5,-78</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-85.5,43,-85.5</points>
<intersection>26.5 0</intersection>
<intersection>43 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>43,-85.5,43,-84.5</points>
<intersection>-85.5 1</intersection>
<intersection>-84.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>43,-84.5,45,-84.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>43 2</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>102,-28,129,-28</points>
<connection>
<GID>150</GID>
<name>CLK</name></connection>
<intersection>103 9</intersection>
<intersection>113 8</intersection>
<intersection>129 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>129,-28,129,-23</points>
<intersection>-28 4</intersection>
<intersection>-23 12</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>113,-28,113,-23</points>
<intersection>-28 4</intersection>
<intersection>-23 11</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>103,-28,103,-23</points>
<intersection>-28 4</intersection>
<intersection>-23 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>103,-23,105,-23</points>
<connection>
<GID>146</GID>
<name>clock</name></connection>
<intersection>103 9</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>113,-23,115,-23</points>
<connection>
<GID>147</GID>
<name>clock</name></connection>
<intersection>113 8</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>129,-23,131,-23</points>
<connection>
<GID>148</GID>
<name>clock</name></connection>
<intersection>129 7</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-25,104,-16</points>
<intersection>-25 4</intersection>
<intersection>-21 3</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>101,-16,104,-16</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104,-21,105,-21</points>
<connection>
<GID>146</GID>
<name>J</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104,-25,105,-25</points>
<connection>
<GID>146</GID>
<name>K</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-21,115,-21</points>
<connection>
<GID>147</GID>
<name>J</name></connection>
<connection>
<GID>146</GID>
<name>Q</name></connection>
<intersection>112 5</intersection>
<intersection>114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114,-25,114,-21</points>
<intersection>-25 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>114,-25,115,-25</points>
<connection>
<GID>147</GID>
<name>K</name></connection>
<intersection>114 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>112,-30,112,-14</points>
<intersection>-30 6</intersection>
<intersection>-21 1</intersection>
<intersection>-14 9</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>112,-30,139,-30</points>
<intersection>112 5</intersection>
<intersection>139 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>139,-30,139,-23</points>
<intersection>-30 6</intersection>
<intersection>-23 11</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>112,-14,123,-14</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>112 5</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>139,-23,140,-23</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>139 7</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-25,130,-15</points>
<intersection>-25 8</intersection>
<intersection>-21 7</intersection>
<intersection>-15 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>129,-15,130,-15</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>130,-21,131,-21</points>
<connection>
<GID>148</GID>
<name>J</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>130,-25,131,-25</points>
<connection>
<GID>148</GID>
<name>K</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-29,122,-16</points>
<intersection>-29 3</intersection>
<intersection>-21 2</intersection>
<intersection>-16 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>121,-21,122,-21</points>
<connection>
<GID>147</GID>
<name>Q</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>122,-29,138,-29</points>
<intersection>122 0</intersection>
<intersection>138 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>138,-29,138,-22</points>
<intersection>-29 3</intersection>
<intersection>-22 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>122,-16,123,-16</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>138,-22,140,-22</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>138 4</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137,-21,140,-21</points>
<connection>
<GID>152</GID>
<name>IN_2</name></connection>
<connection>
<GID>148</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>102,-55,129,-55</points>
<connection>
<GID>158</GID>
<name>CLK</name></connection>
<intersection>103 9</intersection>
<intersection>113 8</intersection>
<intersection>129 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>129,-55,129,-50</points>
<intersection>-55 4</intersection>
<intersection>-50 12</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>113,-55,113,-50</points>
<intersection>-55 4</intersection>
<intersection>-50 11</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>103,-55,103,-50</points>
<intersection>-55 4</intersection>
<intersection>-50 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>103,-50,105,-50</points>
<connection>
<GID>154</GID>
<name>clock</name></connection>
<intersection>103 9</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>113,-50,115,-50</points>
<connection>
<GID>155</GID>
<name>clock</name></connection>
<intersection>113 8</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>129,-50,131,-50</points>
<connection>
<GID>156</GID>
<name>clock</name></connection>
<intersection>129 7</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-52,104,-43</points>
<intersection>-52 4</intersection>
<intersection>-48 3</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>101,-43,104,-43</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104,-48,105,-48</points>
<connection>
<GID>154</GID>
<name>J</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>104,-52,105,-52</points>
<connection>
<GID>154</GID>
<name>K</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-52,130,-42</points>
<intersection>-52 8</intersection>
<intersection>-48 7</intersection>
<intersection>-42 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>129,-42,130,-42</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>130,-48,131,-48</points>
<connection>
<GID>156</GID>
<name>J</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>130,-52,131,-52</points>
<connection>
<GID>156</GID>
<name>K</name></connection>
<intersection>130 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137,-48,140,-48</points>
<connection>
<GID>160</GID>
<name>IN_2</name></connection>
<connection>
<GID>156</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-52,115,-52</points>
<connection>
<GID>155</GID>
<name>K</name></connection>
<connection>
<GID>154</GID>
<name>nQ</name></connection>
<intersection>114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114,-52,114,-41</points>
<intersection>-52 1</intersection>
<intersection>-48 4</intersection>
<intersection>-41 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>114,-48,115,-48</points>
<connection>
<GID>155</GID>
<name>J</name></connection>
<intersection>114 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>114,-41,123,-41</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>114 3</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-52,122,-43</points>
<intersection>-52 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-52,122,-52</points>
<connection>
<GID>155</GID>
<name>nQ</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122,-43,123,-43</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-56,123,-48</points>
<intersection>-56 2</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-48,123,-48</points>
<connection>
<GID>155</GID>
<name>Q</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123,-56,138,-56</points>
<intersection>123 0</intersection>
<intersection>138 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>138,-56,138,-49</points>
<intersection>-56 2</intersection>
<intersection>-49 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>138,-49,140,-49</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>138 3</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>112,-57,139,-57</points>
<intersection>112 4</intersection>
<intersection>139 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>139,-57,139,-50</points>
<intersection>-57 1</intersection>
<intersection>-50 7</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>112,-57,112,-48</points>
<intersection>-57 1</intersection>
<intersection>-48 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>111,-48,112,-48</points>
<connection>
<GID>154</GID>
<name>Q</name></connection>
<intersection>112 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>139,-50,140,-50</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>139 3</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>101,-81.5,146,-81.5</points>
<connection>
<GID>166</GID>
<name>CLK</name></connection>
<intersection>102 9</intersection>
<intersection>113 8</intersection>
<intersection>134 16</intersection>
<intersection>146 15</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>113,-81.5,113,-77</points>
<intersection>-81.5 4</intersection>
<intersection>-77 11</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>102,-81.5,102,-77</points>
<intersection>-81.5 4</intersection>
<intersection>-77 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>102,-77,104,-77</points>
<connection>
<GID>162</GID>
<name>clock</name></connection>
<intersection>102 9</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>113,-77,120,-77</points>
<connection>
<GID>163</GID>
<name>clock</name></connection>
<intersection>113 8</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>146,-81.5,146,-75.5</points>
<intersection>-81.5 4</intersection>
<intersection>-75.5 18</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>134,-81.5,134,-76.5</points>
<intersection>-81.5 4</intersection>
<intersection>-76.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>134,-76.5,136,-76.5</points>
<connection>
<GID>164</GID>
<name>clock</name></connection>
<intersection>134 16</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>146,-75.5,155,-75.5</points>
<connection>
<GID>169</GID>
<name>clock</name></connection>
<intersection>146 15</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-79,103,-70</points>
<intersection>-79 6</intersection>
<intersection>-75 5</intersection>
<intersection>-70 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>101,-70,103,-70</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>103,-75,104,-75</points>
<connection>
<GID>162</GID>
<name>J</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>103,-79,104,-79</points>
<connection>
<GID>162</GID>
<name>K</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>145,-82,163,-82</points>
<intersection>145 6</intersection>
<intersection>163 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>163,-82,163,-74.5</points>
<intersection>-82 1</intersection>
<intersection>-74.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>163,-74.5,166,-74.5</points>
<connection>
<GID>168</GID>
<name>IN_2</name></connection>
<intersection>163 2</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>145,-82,145,-71.5</points>
<intersection>-82 1</intersection>
<intersection>-74.5 7</intersection>
<intersection>-71.5 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>142,-74.5,145,-74.5</points>
<connection>
<GID>164</GID>
<name>Q</name></connection>
<intersection>145 6</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>145,-71.5,147,-71.5</points>
<connection>
<GID>171</GID>
<name>IN_2</name></connection>
<intersection>145 6</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-83,127,-68.5</points>
<intersection>-83 2</intersection>
<intersection>-75 1</intersection>
<intersection>-72 10</intersection>
<intersection>-68.5 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-75,127,-75</points>
<connection>
<GID>163</GID>
<name>Q</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,-83,164,-83</points>
<intersection>127 0</intersection>
<intersection>164 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>164,-83,164,-75.5</points>
<intersection>-83 2</intersection>
<intersection>-75.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>164,-75.5,166,-75.5</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>164 5</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>127,-68.5,128,-68.5</points>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>127,-72,144,-72</points>
<intersection>127 0</intersection>
<intersection>144 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>144,-72,144,-69.5</points>
<intersection>-72 10</intersection>
<intersection>-69.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>144,-69.5,147,-69.5</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>144 11</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161,-73.5,166,-73.5</points>
<connection>
<GID>169</GID>
<name>Q</name></connection>
<connection>
<GID>168</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-64,162,-64</points>
<intersection>111 7</intersection>
<intersection>162 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>162,-77.5,162,-64</points>
<intersection>-77.5 5</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>161,-77.5,162,-77.5</points>
<connection>
<GID>169</GID>
<name>nQ</name></connection>
<intersection>162 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>111,-66.5,111,-64</points>
<intersection>-66.5 8</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>111,-66.5,112,-66.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>111 7</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>112,-84,165,-84</points>
<intersection>112 4</intersection>
<intersection>154 18</intersection>
<intersection>165 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>165,-84,165,-76.5</points>
<intersection>-84 1</intersection>
<intersection>-76.5 13</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>112,-84,112,-70.5</points>
<intersection>-84 1</intersection>
<intersection>-75 5</intersection>
<intersection>-70.5 7</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>110,-75,112,-75</points>
<connection>
<GID>162</GID>
<name>Q</name></connection>
<intersection>112 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>112,-70.5,143,-70.5</points>
<intersection>112 4</intersection>
<intersection>120 10</intersection>
<intersection>125.5 8</intersection>
<intersection>143 16</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>125.5,-70.5,125.5,-66.5</points>
<intersection>-70.5 7</intersection>
<intersection>-66.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>125.5,-66.5,128,-66.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>125.5 8</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>120,-79,120,-70.5</points>
<connection>
<GID>163</GID>
<name>K</name></connection>
<intersection>-70.5 7</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>165,-76.5,166,-76.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>165 3</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>143,-70.5,143,-67.5</points>
<intersection>-70.5 7</intersection>
<intersection>-67.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>143,-67.5,147,-67.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>143 16</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>154,-84,154,-77.5</points>
<intersection>-84 1</intersection>
<intersection>-77.5 19</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>154,-77.5,155,-77.5</points>
<connection>
<GID>169</GID>
<name>K</name></connection>
<intersection>154 18</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-79,111,-68.5</points>
<intersection>-79 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-68.5,112,-68.5</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-79,111,-79</points>
<connection>
<GID>162</GID>
<name>nQ</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-75,119,-67.5</points>
<intersection>-75 1</intersection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-75,120,-75</points>
<connection>
<GID>163</GID>
<name>J</name></connection>
<intersection>119 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118,-67.5,119,-67.5</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-78.5,135,-67.5</points>
<intersection>-78.5 5</intersection>
<intersection>-74.5 3</intersection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>134,-67.5,135,-67.5</points>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>135,-74.5,136,-74.5</points>
<connection>
<GID>164</GID>
<name>J</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>135,-78.5,136,-78.5</points>
<connection>
<GID>164</GID>
<name>K</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-73.5,154,-69.5</points>
<intersection>-73.5 1</intersection>
<intersection>-69.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-73.5,155,-73.5</points>
<connection>
<GID>169</GID>
<name>J</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>153,-69.5,154,-69.5</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>154 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-114.5,151,-114.5</points>
<connection>
<GID>175</GID>
<name>CLK</name></connection>
<intersection>125 14</intersection>
<intersection>141 13</intersection>
<intersection>151 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>151,-114.5,151,-106</points>
<intersection>-114.5 1</intersection>
<intersection>-106 17</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>141,-114.5,141,-106</points>
<intersection>-114.5 1</intersection>
<intersection>-106 16</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>125,-114.5,125,-106</points>
<intersection>-114.5 1</intersection>
<intersection>-106 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>125,-106,127,-106</points>
<connection>
<GID>172</GID>
<name>clock</name></connection>
<intersection>125 14</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>141,-106,143,-106</points>
<connection>
<GID>173</GID>
<name>clock</name></connection>
<intersection>141 13</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>151,-106,153,-106</points>
<connection>
<GID>174</GID>
<name>clock</name></connection>
<intersection>151 12</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-102,119,-100</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>-102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-102,119,-102</points>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119,-98,119,-96</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-96,119,-96</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<intersection>119 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-108,126,-99</points>
<intersection>-108 4</intersection>
<intersection>-104 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-104,127,-104</points>
<connection>
<GID>172</GID>
<name>J</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-99,126,-99</points>
<connection>
<GID>178</GID>
<name>OUT</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>126,-108,127,-108</points>
<connection>
<GID>172</GID>
<name>K</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-111,133.5,-111</points>
<intersection>111 3</intersection>
<intersection>133.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111,-111,111,-103</points>
<intersection>-111 1</intersection>
<intersection>-103 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>133.5,-111,133.5,-108</points>
<intersection>-111 1</intersection>
<intersection>-108 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>111,-103,112,-103</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>111 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>133,-108,133.5,-108</points>
<connection>
<GID>172</GID>
<name>nQ</name></connection>
<intersection>133.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-112,160,-112</points>
<intersection>110 3</intersection>
<intersection>160 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,-112,110,-101</points>
<intersection>-112 1</intersection>
<intersection>-101 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>160,-112,160,-108</points>
<intersection>-112 1</intersection>
<intersection>-108 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>110,-101,112,-101</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>110 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>159,-108,160,-108</points>
<connection>
<GID>174</GID>
<name>nQ</name></connection>
<intersection>160 4</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-93,152,-93</points>
<intersection>111 4</intersection>
<intersection>152 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>152,-116,152,-93</points>
<intersection>-116 8</intersection>
<intersection>-108 11</intersection>
<intersection>-104 16</intersection>
<intersection>-93 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>111,-95,111,-93</points>
<intersection>-95 5</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>111,-95,112,-95</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>111 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>152,-116,162,-116</points>
<intersection>152 3</intersection>
<intersection>162 12</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>152,-108,153,-108</points>
<connection>
<GID>174</GID>
<name>K</name></connection>
<intersection>152 3</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>162,-116,162,-105</points>
<intersection>-116 8</intersection>
<intersection>-105 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>162,-105,164,-105</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>162 12</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>149,-104,153,-104</points>
<connection>
<GID>174</GID>
<name>J</name></connection>
<connection>
<GID>173</GID>
<name>Q</name></connection>
<intersection>152 3</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-92,134,-92</points>
<intersection>110 3</intersection>
<intersection>134 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,-97,110,-92</points>
<intersection>-97 4</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>110,-97,112,-97</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>110 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>134,-117,134,-92</points>
<intersection>-117 6</intersection>
<intersection>-104 11</intersection>
<intersection>-101.5 9</intersection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>134,-117,163,-117</points>
<intersection>134 5</intersection>
<intersection>163 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>163,-117,163,-106</points>
<intersection>-117 6</intersection>
<intersection>-106 10</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>134,-101.5,135.5,-101.5</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>134 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>163,-106,164,-106</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>163 7</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>133,-104,134,-104</points>
<connection>
<GID>172</GID>
<name>Q</name></connection>
<intersection>134 5</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135,-97.5,160,-97.5</points>
<intersection>135 4</intersection>
<intersection>160 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>160,-104,160,-97.5</points>
<intersection>-104 6</intersection>
<intersection>-97.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>135,-99.5,135,-97.5</points>
<intersection>-99.5 7</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>159,-104,164,-104</points>
<connection>
<GID>180</GID>
<name>IN_2</name></connection>
<connection>
<GID>174</GID>
<name>Q</name></connection>
<intersection>160 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>135,-99.5,135.5,-99.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>135 4</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-108,142,-100.5</points>
<intersection>-108 4</intersection>
<intersection>-104 1</intersection>
<intersection>-100.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-104,143,-104</points>
<connection>
<GID>173</GID>
<name>J</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>142,-108,143,-108</points>
<connection>
<GID>173</GID>
<name>K</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>141.5,-100.5,142,-100.5</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>188,-19,192,-19</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<connection>
<GID>215</GID>
<name>OUT_0</name></connection>
<intersection>191 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>191,-25,191,-19</points>
<intersection>-25 10</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>191,-25,200.5,-25</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>191 9</intersection>
<intersection>197 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>197,-25,197,-16</points>
<intersection>-25 10</intersection>
<intersection>-16 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>197,-16,222,-16</points>
<intersection>197 11</intersection>
<intersection>222 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>222,-20,222,-16</points>
<intersection>-20 14</intersection>
<intersection>-16 12</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>222,-20,226,-20</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>222 13</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-33,190,-25</points>
<intersection>-33 4</intersection>
<intersection>-29 1</intersection>
<intersection>-25 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,-29,191,-29</points>
<connection>
<GID>218</GID>
<name>J</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>190,-33,191,-33</points>
<connection>
<GID>218</GID>
<name>K</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>188,-25,190,-25</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>206,-20,207,-20</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<intersection>207 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>207,-22,207,-20</points>
<intersection>-22 7</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>207,-22,208,-22</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>207 3</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-26,207,-24</points>
<intersection>-26 3</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,-24,208,-24</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>206.5,-26,207,-26</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196,-19,200,-19</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>200 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>200,-19,200,-12</points>
<intersection>-19 1</intersection>
<intersection>-12 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>200,-12,226,-12</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>200 5</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-33,198,-14</points>
<intersection>-33 2</intersection>
<intersection>-21 1</intersection>
<intersection>-14 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,-21,200,-21</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-33,198,-33</points>
<connection>
<GID>218</GID>
<name>nQ</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>198,-14,226,-14</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>198 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-35,199,-27</points>
<intersection>-35 4</intersection>
<intersection>-29 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199,-27,200.5,-27</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<intersection>199 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>197,-29,199,-29</points>
<connection>
<GID>218</GID>
<name>Q</name></connection>
<intersection>199 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>199,-35,250,-35</points>
<intersection>199 0</intersection>
<intersection>223 5</intersection>
<intersection>250 7</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>223,-35,223,-22</points>
<intersection>-35 4</intersection>
<intersection>-22 9</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>250,-35,250,-29</points>
<intersection>-35 4</intersection>
<intersection>-29 10</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>223,-22,226,-22</points>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<intersection>223 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>250,-29,251,-29</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>250 7</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>215,-31,215,-23</points>
<intersection>-31 4</intersection>
<intersection>-27 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>215,-27,216,-27</points>
<connection>
<GID>219</GID>
<name>J</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214,-23,215,-23</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<intersection>215 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>215,-31,216,-31</points>
<connection>
<GID>219</GID>
<name>K</name></connection>
<intersection>215 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-31,225,-16</points>
<intersection>-31 2</intersection>
<intersection>-16 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>222,-31,225,-31</points>
<connection>
<GID>219</GID>
<name>nQ</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>225,-16,226,-16</points>
<connection>
<GID>209</GID>
<name>IN_2</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>224,-34,224,-24</points>
<intersection>-34 1</intersection>
<intersection>-27 2</intersection>
<intersection>-24 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>224,-34,249,-34</points>
<intersection>224 0</intersection>
<intersection>249 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>222,-27,224,-27</points>
<connection>
<GID>219</GID>
<name>Q</name></connection>
<intersection>224 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>249,-34,249,-28</points>
<intersection>-34 1</intersection>
<intersection>-28 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>249,-28,251,-28</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>249 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>224,-24,226,-24</points>
<connection>
<GID>210</GID>
<name>IN_2</name></connection>
<intersection>224 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-17,233,-14</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-14 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>232,-14,233,-14</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<intersection>233 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>233,-22,233,-19</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>-22 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>232,-22,233,-22</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<intersection>233 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>240,-31,240,-18</points>
<intersection>-31 4</intersection>
<intersection>-27 1</intersection>
<intersection>-18 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>240,-27,241,-27</points>
<connection>
<GID>220</GID>
<name>J</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>240,-31,241,-31</points>
<connection>
<GID>220</GID>
<name>K</name></connection>
<intersection>240 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>239,-18,240,-18</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>240 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>247,-27,251,-27</points>
<connection>
<GID>220</GID>
<name>Q</name></connection>
<connection>
<GID>212</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>188,-38,239,-38</points>
<connection>
<GID>213</GID>
<name>CLK</name></connection>
<intersection>189 4</intersection>
<intersection>214 9</intersection>
<intersection>239 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>189,-38,189,-31</points>
<intersection>-38 1</intersection>
<intersection>-31 12</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>239,-38,239,-29</points>
<intersection>-38 1</intersection>
<intersection>-29 11</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>214,-38,214,-29</points>
<intersection>-38 1</intersection>
<intersection>-29 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>214,-29,216,-29</points>
<connection>
<GID>219</GID>
<name>clock</name></connection>
<intersection>214 9</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>239,-29,241,-29</points>
<connection>
<GID>220</GID>
<name>clock</name></connection>
<intersection>239 8</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>189,-31,191,-31</points>
<connection>
<GID>218</GID>
<name>clock</name></connection>
<intersection>189 4</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>20.925,-0.790047,211.587,-95.0304</PageViewport>
<gate>
<ID>238</ID>
<type>AA_LABEL</type>
<position>60,-63.5</position>
<gparam>LABEL_TEXT Ring Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>239</ID>
<type>AE_DFF_LOW</type>
<position>46,-75.5</position>
<input>
<ID>IN_0</ID>201 </input>
<output>
<ID>OUT_0</ID>197 </output>
<input>
<ID>clock</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>240</ID>
<type>AE_DFF_LOW</type>
<position>57,-75.5</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>198 </output>
<input>
<ID>clock</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_DFF_LOW</type>
<position>68,-75.5</position>
<input>
<ID>IN_0</ID>198 </input>
<output>
<ID>OUT_0</ID>199 </output>
<input>
<ID>clock</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>242</ID>
<type>AE_DFF_LOW</type>
<position>79,-75.5</position>
<input>
<ID>IN_0</ID>199 </input>
<output>
<ID>OUT_0</ID>201 </output>
<input>
<ID>clock</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>243</ID>
<type>BB_CLOCK</type>
<position>37,-83.5</position>
<output>
<ID>CLK</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>244</ID>
<type>GA_LED</type>
<position>51,-70.5</position>
<input>
<ID>N_in2</ID>197 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>GA_LED</type>
<position>63,-70.5</position>
<input>
<ID>N_in2</ID>198 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>GA_LED</type>
<position>73.5,-70.5</position>
<input>
<ID>N_in2</ID>199 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>GA_LED</type>
<position>85,-70.5</position>
<input>
<ID>N_in2</ID>201 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,-73.5,54,-73.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<connection>
<GID>239</GID>
<name>OUT_0</name></connection>
<intersection>51 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51,-73.5,51,-71.5</points>
<connection>
<GID>244</GID>
<name>N_in2</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-73.5,65,-73.5</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>63 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-73.5,63,-71.5</points>
<connection>
<GID>245</GID>
<name>N_in2</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,-73.5,76,-73.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<intersection>73.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73.5,-73.5,73.5,-71.5</points>
<connection>
<GID>246</GID>
<name>N_in2</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41,-83.5,75,-83.5</points>
<connection>
<GID>243</GID>
<name>CLK</name></connection>
<intersection>42 9</intersection>
<intersection>53 8</intersection>
<intersection>64 7</intersection>
<intersection>75 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>75,-83.5,75,-76.5</points>
<intersection>-83.5 1</intersection>
<intersection>-76.5 13</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>64,-83.5,64,-76.5</points>
<intersection>-83.5 1</intersection>
<intersection>-76.5 11</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>53,-83.5,53,-76.5</points>
<intersection>-83.5 1</intersection>
<intersection>-76.5 12</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>42,-83.5,42,-76.5</points>
<intersection>-83.5 1</intersection>
<intersection>-76.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>42,-76.5,43,-76.5</points>
<connection>
<GID>239</GID>
<name>clock</name></connection>
<intersection>42 9</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>64,-76.5,65,-76.5</points>
<connection>
<GID>241</GID>
<name>clock</name></connection>
<intersection>64 7</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>53,-76.5,54,-76.5</points>
<connection>
<GID>240</GID>
<name>clock</name></connection>
<intersection>53 8</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>75,-76.5,76,-76.5</points>
<connection>
<GID>242</GID>
<name>clock</name></connection>
<intersection>75 6</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-68.5,83,-68.5</points>
<intersection>42 5</intersection>
<intersection>83 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>83,-73.5,83,-68.5</points>
<intersection>-73.5 8</intersection>
<intersection>-68.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>42,-73.5,42,-68.5</points>
<intersection>-73.5 10</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>82,-73.5,85,-73.5</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>83 4</intersection>
<intersection>85 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>85,-73.5,85,-71.5</points>
<connection>
<GID>247</GID>
<name>N_in2</name></connection>
<intersection>-73.5 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>42,-73.5,43,-73.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>42 5</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>42.3692,12.6731,296.585,-112.981</PageViewport>
<gate>
<ID>260</ID>
<type>AA_LABEL</type>
<position>48,-16</position>
<gparam>LABEL_TEXT Twisted Ring Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>AE_DFF_LOW</type>
<position>32,-28.5</position>
<input>
<ID>IN_0</ID>213 </input>
<output>
<ID>OUT_0</ID>209 </output>
<input>
<ID>clock</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>262</ID>
<type>AE_DFF_LOW</type>
<position>43,-28.5</position>
<input>
<ID>IN_0</ID>209 </input>
<output>
<ID>OUT_0</ID>210 </output>
<input>
<ID>clock</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>263</ID>
<type>AE_DFF_LOW</type>
<position>54,-28.5</position>
<input>
<ID>IN_0</ID>210 </input>
<output>
<ID>OUT_0</ID>211 </output>
<input>
<ID>clock</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>264</ID>
<type>AE_DFF_LOW</type>
<position>65,-28.5</position>
<input>
<ID>IN_0</ID>211 </input>
<output>
<ID>OUTINV_0</ID>213 </output>
<output>
<ID>OUT_0</ID>214 </output>
<input>
<ID>clock</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>265</ID>
<type>BB_CLOCK</type>
<position>23,-36.5</position>
<output>
<ID>CLK</ID>212 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>266</ID>
<type>GA_LED</type>
<position>37,-23.5</position>
<input>
<ID>N_in2</ID>209 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>GA_LED</type>
<position>49,-23.5</position>
<input>
<ID>N_in2</ID>210 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>GA_LED</type>
<position>59.5,-23.5</position>
<input>
<ID>N_in2</ID>211 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>GA_LED</type>
<position>71,-23.5</position>
<input>
<ID>N_in2</ID>214 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-26.5,40,-26.5</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>37 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37,-26.5,37,-24.5</points>
<connection>
<GID>266</GID>
<name>N_in2</name></connection>
<intersection>-26.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46,-26.5,51,-26.5</points>
<connection>
<GID>262</GID>
<name>OUT_0</name></connection>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>49 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49,-26.5,49,-24.5</points>
<connection>
<GID>267</GID>
<name>N_in2</name></connection>
<intersection>-26.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-26.5,62,-26.5</points>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>59.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>59.5,-26.5,59.5,-24.5</points>
<connection>
<GID>268</GID>
<name>N_in2</name></connection>
<intersection>-26.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-36.5,61,-36.5</points>
<connection>
<GID>265</GID>
<name>CLK</name></connection>
<intersection>28 9</intersection>
<intersection>39 8</intersection>
<intersection>50 7</intersection>
<intersection>61 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>61,-36.5,61,-29.5</points>
<intersection>-36.5 1</intersection>
<intersection>-29.5 13</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>50,-36.5,50,-29.5</points>
<intersection>-36.5 1</intersection>
<intersection>-29.5 11</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>39,-36.5,39,-29.5</points>
<intersection>-36.5 1</intersection>
<intersection>-29.5 12</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>28,-36.5,28,-29.5</points>
<intersection>-36.5 1</intersection>
<intersection>-29.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>28,-29.5,29,-29.5</points>
<connection>
<GID>261</GID>
<name>clock</name></connection>
<intersection>28 9</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>50,-29.5,51,-29.5</points>
<connection>
<GID>263</GID>
<name>clock</name></connection>
<intersection>50 7</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>39,-29.5,40,-29.5</points>
<connection>
<GID>262</GID>
<name>clock</name></connection>
<intersection>39 8</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>61,-29.5,62,-29.5</points>
<connection>
<GID>264</GID>
<name>clock</name></connection>
<intersection>61 6</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-20.5,69,-20.5</points>
<intersection>28 3</intersection>
<intersection>69 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28,-26.5,28,-20.5</points>
<intersection>-26.5 4</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>28,-26.5,29,-26.5</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>28 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>69,-29.5,69,-20.5</points>
<intersection>-29.5 6</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>68,-29.5,69,-29.5</points>
<connection>
<GID>264</GID>
<name>OUTINV_0</name></connection>
<intersection>69 5</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-26.5,71,-24.5</points>
<connection>
<GID>269</GID>
<name>N_in2</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-26.5,71,-26.5</points>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 3>
<page 4>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 4>
<page 5>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 5>
<page 6>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 6>
<page 7>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 7>
<page 8>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 8>
<page 9>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 9></circuit>